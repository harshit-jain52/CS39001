`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.09.2024 16:08:49
// Design Name: 
// Module Name: multN
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module multN #(parameter N = 8)(
    input wire [N-1:0] A, B,
    output wire [N-1:0] P
    );
    
    assign P = A * B;
endmodule
