module ins_mem(
    input wire rst,
	input [31:0] addr,
	output reg [31:0] ins
);
	reg [31:0] mem [1023:0];
	
//	initial begin
//		$readmemb("sum10_ins_bin.mem", mem, 0, 1023);
//		$monitor("Time:%0t | PC = %d, ins = %b", $time, addr[9:0], mem[addr[9:0]]);
//	end
    
    always@(posedge rst) begin
        // Sum of natural numbers till 10
//        mem[0] <= 32'b01000100000000010000000000000000;
//        mem[1] <= 32'b10001100001000000000000000000100;
//        mem[2] <= 32'b00000000010000010001000000000001;
//        mem[3] <= 32'b00001000001000010000000000000001;
//        mem[4] <= 32'b10000011111111111111111111111101;
//        mem[5] <= 32'b10010000000000000000000000000000;

        // Insertion sort of 10 integers 
        mem[0] <= 32'b00000100000000010000000000000001;
        mem[1] <= 32'b00101000001001000000000000001010;
        mem[2] <= 32'b10001100100000000000000000001101;
        mem[3] <= 32'b00001000001000100000000000000001;
        mem[4] <= 32'b01000100001000110000000000000000;
        mem[5] <= 32'b10000100010000000000000000000111;
        mem[6] <= 32'b01000100010001010000000000000000;
        mem[7] <= 32'b00000000011001010010000000001010;
        mem[8] <= 32'b10001100100000000000000000000100;
        mem[9] <= 32'b01001000010001010000000000000001;
        mem[10] <= 32'b00000000000000100001000000001110;
        mem[11] <= 32'b10000011111111111111111111111010;
        mem[12] <= 32'b01001000010000110000000000000001;
        mem[13] <= 32'b00000000000000010000100000001101;
        mem[14] <= 32'b10000011111111111111111111110011;
        mem[15] <= 32'b01000100000000010000000000000000;
        mem[16] <= 32'b01000100000000100000000000000001;
        mem[17] <= 32'b01000100000000110000000000000010;
        mem[18] <= 32'b01000100000001000000000000000011;
        mem[19] <= 32'b01000100000001010000000000000100;
        mem[20] <= 32'b01000100000001100000000000000101;
        mem[21] <= 32'b01000100000001110000000000000110;
        mem[22] <= 32'b01000100000010000000000000000111;
        mem[23] <= 32'b01000100000010010000000000001000;
        mem[24] <= 32'b01000100000010100000000000001001;
        mem[25] <= 32'b10010000000000000000000000000000;
    end
    
	always @(*) begin 
//		 $display("PC = %d, ins = %b", addr[9:0], mem[addr[9:0]]);
		ins = mem[addr[9:0]];
	end
endmodule