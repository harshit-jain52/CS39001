module mux16x1N_tb;
    parameter N = 8; 
    reg [N-1:0] D [15:0]; 
    reg [3:0] S;           
    wire [N-1:0] Z;       
    
    mux16x1N #(N) uut (.D(D), .S(S), .Z(Z));

    initial begin
        $monitor("Time = %0t | S = %b | Z = %d", $time, S, Z);

        D[0] = 8'b0000_0001;
        D[1] = 8'b0000_0010;
        D[2] = 8'b0000_0100;
        D[3] = 8'b0000_1000;
        D[4] = 8'b0001_0000;
        D[5] = 8'b0010_0000;
        D[6] = 8'b0100_0000;
        D[7] = 8'b1000_0000;
        D[8] = 8'b1111_0000;
        D[9] = 8'b1110_0000;
        D[10] = 8'b1100_0000;
        D[11] = 8'b1000_0000;
        D[12] = 8'b0000_1111;
        D[13] = 8'b0000_1110;
        D[14] = 8'b0000_1100;
        D[15] = 8'b0000_1000;

        $display("D = %p", D);

        S = 4'b0000; #10; 
        S = 4'b0001; #10; 
        S = 4'b0010; #10; 
        S = 4'b0011; #10; 
        S = 4'b0100; #10; 
        S = 4'b0101; #10; 
        S = 4'b0110; #10; 
        S = 4'b0111; #10; 
        S = 4'b1000; #10; 
        S = 4'b1001; #10; 
        S = 4'b1010; #10; 
        S = 4'b1011; #10; 
        S = 4'b1100; #10; 
        S = 4'b1101; #10; 
        S = 4'b1110; #10; 
        S = 4'b1111; #10; 

        #100 $finish;
    end

endmodule
